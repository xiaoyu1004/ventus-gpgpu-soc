`timescale 1ns/10ps

`include "define.v"

module gpgpu_top_wrapper (
  input clk,
  input rst_n,

  input                           host_req_valid_i,
  output                          host_req_ready_o,
  input  [      `WG_ID_WIDTH-1:0] host_req_wg_id_i,
  input  [   `WF_COUNT_WIDTH-1:0] host_req_num_wf_i,
  input  [  `WAVE_ITEM_WIDTH-1:0] host_req_wf_size_i,
  input  [   `MEM_ADDR_WIDTH-1:0] host_req_start_pc_i,
  input  [`WG_SIZE_X_WIDTH-1:0]   host_req_kernel_size_x_i,
  input  [`WG_SIZE_X_WIDTH-1:0]   host_req_kernel_size_y_i,
  input  [`WG_SIZE_X_WIDTH-1:0]   host_req_kernel_size_z_i,
  input  [   `MEM_ADDR_WIDTH-1:0] host_req_pds_baseaddr_i,
  input  [   `MEM_ADDR_WIDTH-1:0] host_req_csr_knl_i,
  input  [      `VGPR_ID_WIDTH:0] host_req_vgpr_size_total_i,
  input  [      `SGPR_ID_WIDTH:0] host_req_sgpr_size_total_i,
  input  [       `LDS_ID_WIDTH:0] host_req_lds_size_total_i,
  input  [       `GDS_ID_WIDTH:0] host_req_gds_size_total_i,
  input  [      `VGPR_ID_WIDTH:0] host_req_vgpr_size_per_wf_i,
  input  [      `SGPR_ID_WIDTH:0] host_req_sgpr_size_per_wf_i,
  input  [   `MEM_ADDR_WIDTH-1:0] host_req_gds_baseaddr_i,

  output                    host_rsp_valid_o,
  input                     host_rsp_ready_i,
  output [`WG_ID_WIDTH-1:0] host_rsp_inflight_wg_buffer_host_wf_done_wg_id_o,

  //AXI
  output [                          `NUM_L2CACHE-1:0] out_a_valid_o,
  input  [                          `NUM_L2CACHE-1:0] out_a_ready_i,
  output [                 `NUM_L2CACHE*`OP_BITS-1:0] out_a_opcode_o,
  output [               `NUM_L2CACHE*`SIZE_BITS-1:0] out_a_size_o,
  output [             `NUM_L2CACHE*`SOURCE_BITS-1:0] out_a_source_o,
  output [            `NUM_L2CACHE*`ADDRESS_BITS-1:0] out_a_address_o,
  output [               `NUM_L2CACHE*`MASK_BITS-1:0] out_a_mask_o,
  output [               `NUM_L2CACHE*`DATA_BITS-1:0] out_a_data_o,
  output [                        `NUM_L2CACHE*3-1:0] out_a_param_o,

  input  [             `NUM_L2CACHE-1:0] out_d_valid_i,
  output [             `NUM_L2CACHE-1:0] out_d_ready_o,
  input  [    `NUM_L2CACHE*`OP_BITS-1:0] out_d_opcode_i,
  input  [  `NUM_L2CACHE*`SIZE_BITS-1:0] out_d_size_i,
  input  [`NUM_L2CACHE*`SOURCE_BITS-1:0] out_d_source_i,
  input  [  `NUM_L2CACHE*`DATA_BITS-1:0] out_d_data_i,
  input  [           `NUM_L2CACHE*3-1:0] out_d_param_i
);
  wire [`WG_SIZE_X_WIDTH-1:0]           host_req_kernel_size_3d_i = {host_req_kernel_size_z_i, host_req_kernel_size_y_i, host_req_kernel_size_x_i};

  GPGPU_top gpu_top(
    .clk                                              (clk                                             ),
    .rst_n                                            (rst_n                                           ),
    .host_req_valid_i                                 (host_req_valid_i                                ),
    .host_req_ready_o                                 (host_req_ready_o                                ),
    .host_req_wg_id_i                                 (host_req_wg_id_i                                ),
    .host_req_num_wf_i                                (host_req_num_wf_i                               ),
    .host_req_wf_size_i                               (host_req_wf_size_i                              ),
    .host_req_start_pc_i                              (host_req_start_pc_i                             ),
    .host_req_kernel_size_3d_i                        (host_req_kernel_size_3d_i                       ),
    .host_req_pds_baseaddr_i                          (host_req_pds_baseaddr_i                         ),
    .host_req_csr_knl_i                               (host_req_csr_knl_i                              ),
    .host_req_vgpr_size_total_i                       (host_req_vgpr_size_total_i                      ),
    .host_req_sgpr_size_total_i                       (host_req_sgpr_size_total_i                      ),
    .host_req_lds_size_total_i                        (host_req_lds_size_total_i                       ),
    .host_req_gds_size_total_i                        (host_req_gds_size_total_i                       ),
    .host_req_vgpr_size_per_wf_i                      (host_req_vgpr_size_per_wf_i                     ),
    .host_req_sgpr_size_per_wf_i                      (host_req_sgpr_size_per_wf_i                     ),
    .host_req_gds_baseaddr_i                          (host_req_gds_baseaddr_i                         ),
    .host_rsp_valid_o                                 (host_rsp_valid_o                                ),
    .host_rsp_ready_i                                 (host_rsp_ready_i                                ),
    .host_rsp_inflight_wg_buffer_host_wf_done_wg_id_o (host_rsp_inflight_wg_buffer_host_wf_done_wg_id_o),
    .out_a_valid_o                                    (out_a_valid_o                                   ),
    .out_a_ready_i                                    (out_a_ready_i                                   ),
    .out_a_opcode_o                                   (out_a_opcode_o                                  ),
    .out_a_size_o                                     (out_a_size_o                                    ),
    .out_a_source_o                                   (out_a_source_o                                  ),
    .out_a_address_o                                  (out_a_address_o                                 ),
    .out_a_mask_o                                     (out_a_mask_o                                    ),
    .out_a_data_o                                     (out_a_data_o                                    ),
    .out_a_param_o                                    (out_a_param_o                                   ),
    .out_d_valid_i                                    (out_d_valid_i                                   ),
    .out_d_ready_o                                    (out_d_ready_o                                   ),
    .out_d_opcode_i                                   (out_d_opcode_i                                  ),
    .out_d_size_i                                     (out_d_size_i                                    ),
    .out_d_source_i                                   (out_d_source_i                                  ),
    .out_d_data_i                                     (out_d_data_i                                    ),
    .out_d_param_i                                    (out_d_param_i                                   )
  );

endmodule